--library IEEE;
--use IEEE.STD_LOGIC_1164.ALL;
--
--entity RF_top is
--   port ( 
--
--	);
--end RF_top;
--
--architecture behavioral of RF_top is
--begin
--
--
--end behavioral;